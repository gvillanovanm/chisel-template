module BB (
	input [31:0] io_input,
	output [31:0] io_output
);

assign io_output = io_input;

endmodule